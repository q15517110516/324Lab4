-- ----------------------------------------------------------------------------------
-- -- Company: 
-- -- Engineer: 
-- -- 
-- -- Create Date: 2019/05/09 11:18:41
-- -- Design Name: 
-- -- Module Name: MUX - Behavioral
-- -- Project Name: 
-- -- Target Devices: 
-- -- Tool Versions: 
-- -- Description: 
-- -- 
-- -- Dependencies: 
-- -- 
-- -- Revision:
-- -- Revision 0.01 - File Created
-- -- Additional Comments:
-- -- 
-- ----------------------------------------------------------------------------------


-- LIBRARY IEEE;
-- USE IEEE.STD_LOGIC_1164.ALL;
-- USE IEEE.STD_LOGIC_ARITH.ALL;
-- USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- ENTITY MUX IS
  -- PORT(    
  -- D0       : IN STD_LOGIC_VECTOR(7 DOWNTO 0);--
   -- D1        : IN STD_LOGIC_VECTOR(7 DOWNTO 0);--    
   -- Y        : OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);--
   -- SEL     : IN  STD_LOGIC
      -- );
-- END ENTITY MUX;

-- ARCHITECTURE BEHAV OF MUX IS
-- BEGIN
    
         -- Y <= D0 when SEL='1' else  
              -- D1;    

 -- END ARCHITECTURE BEHAV;